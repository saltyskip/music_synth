module exponential_rom(
		input clk,
		input [5:0] duration,
		output reg [9:0] dout
	);
	wire [9:0] memory [127:0];
	always @(posedge clk)
		dout = memory[duration];
assign memory [0] = {10'd0384};
assign memory [1] = {10'd0512};
assign memory [2] = {10'd0640};
assign memory [3] = {10'd0768};
assign memory [4] = {10'd0896};
assign memory[5] = {10'd1023};
assign memory[6] = {10'd1001};
assign memory[7] = {10'd0981};
assign memory[8] = {10'd0961};
assign memory[9] = {10'd0941};
assign memory[10] = {10'd0921};
assign memory[11] = {10'd0902};
assign memory[12] = {10'd0884};
assign memory[13] = {10'd0865};
assign memory[14] = {10'd0848};
assign memory[15] = {10'd0830};
assign memory[16] = {10'd0813};
assign memory[17] = {10'd0796};
assign memory[18] = {10'd0780};
assign memory[19] = {10'd0764};
assign memory[20] = {10'd0748};
assign memory[21] = {10'd0733};
assign memory[22] = {10'd0717};
assign memory[23] = {10'd0703};
assign memory[24] = {10'd0688};
assign memory[25] = {10'd0674};
assign memory[26] = {10'd0660};
assign memory[27] = {10'd0646};
assign memory[28] = {10'd0633};
assign memory[29] = {10'd0620};
assign memory[30] = {10'd0607};
assign memory[31] = {10'd0595};
assign memory[32] = {10'd0582};
assign memory[33] = {10'd0570};
assign memory[34] = {10'd0559};
assign memory[35] = {10'd0547};
assign memory[36] = {10'd0536};
assign memory[37] = {10'd0525};
assign memory[38] = {10'd0514};
assign memory[39] = {10'd0503};
assign memory[40] = {10'd0493};
assign memory[41] = {10'd0483};
assign memory[42] = {10'd0473};
assign memory[43] = {10'd0463};
assign memory[44] = {10'd0453};
assign memory[45] = {10'd0444};
assign memory[46] = {10'd0435};
assign memory[47] = {10'd0426};
assign memory[48] = {10'd0417};
assign memory[49] = {10'd0409};
assign memory[50] = {10'd0400};
assign memory[51] = {10'd0392};
assign memory[52] = {10'd0384};
assign memory[53] = {10'd0376};
assign memory[54] = {10'd0368};
assign memory[55] = {10'd0360};
assign memory[56] = {10'd0353};
assign memory[57] = {10'd0346};
assign memory[58] = {10'd0339};
assign memory[59] = {10'd0332};
assign memory[60] = {10'd0325};
assign memory[61] = {10'd0318};
assign memory[62] = {10'd0311};
assign memory[63] = {10'd0305};
assign memory[64] = {10'd0299};
assign memory[65] = {10'd0293};
assign memory[66] = {10'd0287};
assign memory[67] = {10'd0281};
assign memory[68] = {10'd0275};
assign memory[69] = {10'd0269};
assign memory[70] = {10'd0264};
assign memory[71] = {10'd0258};
assign memory[72] = {10'd0253};
assign memory[73] = {10'd0248};
assign memory[74] = {10'd0242};
assign memory[75] = {10'd0237};
assign memory[76] = {10'd0233};
assign memory[77] = {10'd0228};
assign memory[78] = {10'd0223};
assign memory[79] = {10'd0218};
assign memory[80] = {10'd0214};
assign memory[81] = {10'd0210};
assign memory[82] = {10'd0205};
assign memory[83] = {10'd0201};
assign memory[84] = {10'd0197};
assign memory[85] = {10'd0193};
assign memory[86] = {10'd0189};
assign memory[87] = {10'd0185};
assign memory[88] = {10'd0181};
assign memory[89] = {10'd0177};
assign memory[90] = {10'd0174};
assign memory[91] = {10'd0170};
assign memory[92] = {10'd0167};
assign memory[93] = {10'd0163};
assign memory[94] = {10'd0160};
assign memory[95] = {10'd0156};
assign memory[96] = {10'd0153};
assign memory[97] = {10'd0150};
assign memory[98] = {10'd0147};
assign memory[99] = {10'd0144};
assign memory[100] = {10'd0141};
assign memory[101] = {10'd0138};
assign memory[102] = {10'd0135};
assign memory[103] = {10'd0132};
assign memory[104] = {10'd0130};
assign memory[105] = {10'd0127};
assign memory[106] = {10'd0124};
assign memory[107] = {10'd0122};
assign memory[108] = {10'd0119};
assign memory[109] = {10'd0117};
assign memory[110] = {10'd0114};
assign memory[111] = {10'd0112};
assign memory[112] = {10'd0110};
assign memory[113] = {10'd0107};
assign memory[114] = {10'd0105};
assign memory[115] = {10'd0103};
assign memory[116] = {10'd0101};
assign memory[117] = {10'd0099};
assign memory[118] = {10'd0097};
assign memory[119] = {10'd0095};
assign memory[120] = {10'd0093};
assign memory[121] = {10'd0091};
assign memory[122] = {10'd0089};
assign memory[123] = {10'd0087};
assign memory[124] = {10'd0085};
assign memory[125] = {10'd0083};
assign memory[126] = {10'd0082};
assign memory[127] = {10'd0080};
endmodule
