//  How to use: 
//  1. Edit the songs on the Enter Song sheet.  
//  2. Select this whole worksheet, copy it, and paste it into a new file.  
//  3. Save the file as song_rom.v. 

module song_rom (
    input clk,
    input [8:0] addr,
    output reg [15:0] dout
);  

    wire [15:0] memory [511:0];

    always @(posedge clk)                       
        dout = memory[addr];                    

    assign memory[   0  ] = {1'b0, 6'd3, 6'd12, 3'b101}  ;   // B       // Lines here test meta=1 (harmonics)
    assign memory[   1  ] = {1'b0, 6'd11, 6'd24, 3'b100}   ;   // G
    assign memory[   2  ] = {1'b0, 6'd18, 6'd12, 3'b100}   ;   // D
    assign memory[   3  ] = {1'b0, 6'd45, 6'd12, 3'b100}   ;   // Note: F
    assign memory[   4  ] = {1'b0, 6'd35, 6'd24, 3'b100}  ;   // Note: G      // G7 chord
    assign memory[   5  ] = {1'b1, 6'd0, 6'd12, 3'b0}  ;   // Note: Advance
    assign memory[   6  ] = {1'b0, 6'd44, 6'd12, 3'b100}  ;   // Note: E
    assign memory[   7  ] = {1'b0, 6'd16, 6'd12, 3'b100}  ;   // Note: C      // resolution to C chord
    assign memory[   8  ] = {1'b1, 6'd0, 6'd12, 3'b0}  ;   // Note: Advance  // end  
    assign memory[   9  ] = {1'b0, 6'd4, 6'd48, 3'b100}   ;   // Note: 1A
    assign memory[   10  ] = {1'b1, 6'd0, 6'd48, 3'b0}   ;   // Advance
    assign memory[   11  ] = {1'b0, 6'd3, 6'd24, 3'b101}   ;   // Note: 1B
    assign memory[   12  ] = {1'b0, 6'd11, 6'd48, 3'b1}  ;   // Note: 1G
    assign memory[   13  ] = {1'b0, 6'd18, 6'd24, 3'b1}  ;   // Note: 2D
    assign memory[   14  ] = {1'b1, 6'd0, 6'd48, 3'b0}   ;   // Advance
    assign memory[   15  ] = {1'b0, 6'd0, 6'd48, 3'b0}   ;   // Rest
    assign memory[   16  ] = {1'b1, 6'd0, 6'd48, 3'b0}  ;  
    assign memory[   17  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   18  ] = {1'b0, 6'd18, 6'd63,3'b110}  ;
    assign memory[   19  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   20  ] = {1'b0, 6'd18, 6'd63,3'b110}  ;
    assign memory[   21  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   22  ] = {1'b0, 6'd18, 6'd63,3'b100}  ;
    assign memory[   23  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   24  ] = {1'b0, 6'd18, 6'd63,3'b100}  ;
    assign memory[   25  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   26  ] = {1'b0, 6'd18, 6'd63,3'b000}  ;
    assign memory[   27  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   28  ] = {1'b0, 6'd18, 6'd63,3'b000}  ;
    assign memory[   29  ] = {1'b1, 6'd0, 6'd63, 3'b0}  ;
    assign memory[   30  ] = {1'b0, 6'd0, 6'd48, 3'b0}  ;  // rest
    assign memory[   31  ] = {1'b1, 6'd0, 6'd48, 3'b0}  ;
    assign memory[   32  ] = {1'b0, 6'd42, 6'd32, 3'b0}  ;  // D
    assign memory[   33  ] = {1'b0, 6'd37, 6'd32, 3'b0}  ;  // A
    assign memory[   34  ] = {1'b0, 6'd33, 6'd32, 3'b0}  ;  // F
    assign memory[   35  ] = {1'b0, 6'd30, 6'd16, 3'b0}  ;  // D
    assign memory[   36  ] = {1'b1, 6'd0, 6'd16, 3'b0}  ;
    assign memory[   37  ] = {1'b0, 6'd18, 6'd16, 3'b0}  ;
    assign memory[   38  ] = {1'b1, 6'd0, 6'd16, 3'b0}  ;
    assign memory[   39  ] = {1'b0, 6'd40, 6'd16, 3'b0}  ;
    assign memory[   40  ] = {1'b0, 6'd35, 6'd16, 3'b0}  ;
    assign memory[   41  ] = {1'b0, 6'd32, 6'd16, 3'b0}  ;
    assign memory[   42  ] = {1'b0, 6'd20, 6'd16, 3'b0}  ;
    assign memory[   43  ] = {1'b1, 6'd0, 6'd16, 3'b0}  ;
    assign memory[   44  ] = {1'b0, 6'd42, 6'd8, 3'b0}  ;
    assign memory[   45  ] = {1'b0, 6'd37, 6'd16, 3'b0}  ;
    assign memory[   46  ] = {1'b0, 6'd30, 6'd32, 3'b0}  ;
    assign memory[   47  ] = {1'b0, 6'd21, 6'd16, 3'b0}  ;
    assign memory[   48  ] = {1'b1, 6'd0, 6'd8, 3'b0}  ;
    assign memory[   49  ] = {1'b0, 6'd40, 6'd8, 3'b0}  ;
    assign memory[   50  ] = {1'b1, 6'd0, 6'd8, 3'b0}  ;
    assign memory[   51  ] = {1'b0, 6'd38, 6'd16, 3'b0}  ;  // Bb
    assign memory[   52  ] = {1'b0, 6'd35, 6'd8, 3'b0}  ;
    assign memory[   53  ] = {1'b0, 6'd23, 6'd16, 3'b0}  ;
    assign memory[   54  ] = {1'b1, 6'd0, 6'd8, 3'b0}  ;
    assign memory[   55  ] = {1'b0, 6'd33, 6'd8, 3'b0}  ;
    assign memory[   56  ] = {1'b1, 6'd0, 6'd8, 3'b0}  ;
    assign memory[   57  ] = {1'b0, 6'd37, 6'd8, 3'b0}  ;
    assign memory[   58  ] = {1'b0, 6'd32, 6'd16, 3'b0}  ;
    assign memory[   59  ] = {1'b0, 6'd29, 6'd16, 3'b0}  ;
    assign memory[   60  ] = {1'b0, 6'd25, 6'd16, 3'b0}  ;
    assign memory[   61  ] = {1'b1, 6'd0, 6'd8, 3'b0}  ;
    assign memory[   62  ] = {1'b0, 6'd35, 6'd8, 3'b0}  ;
    assign memory[   63  ] = {1'b1, 6'd0, 6'd8, 3'b0}  ;
    assign memory[   64  ] = {1'b0, 6'd33, 6'd32, 3'b0}  ;
    assign memory[   65  ] = {1'b0, 6'd30, 6'd48, 3'b0}  ;
    assign memory[   66  ] = {1'b0, 6'd26, 6'd48, 3'b0}  ;
    assign memory[   67  ] = {1'b1, 6'd0, 6'd32, 3'b0}  ;
    assign memory[   68  ] = {1'b0, 6'd35, 6'd16, 3'b0}  ;
    assign memory[   69  ] = {1'b1, 6'd0, 6'd16, 3'b0}  ;
    assign memory[   70  ] = {1'b0, 6'd37, 6'd48, 3'b0}  ;
    assign memory[   71  ] = {1'b0, 6'd32, 6'd48, 3'b0}  ;
    assign memory[   72  ] = {1'b0, 6'd29, 6'd48, 3'b0}  ;
    assign memory[   73  ] = {1'b0, 6'd25, 6'd48, 3'b0}  ;
    assign memory[   74  ] = {1'b1, 6'd0, 6'd48, 3'b0}  ;
    assign memory[   75  ] = {16'b0}  ;
    assign memory[   76  ] = {16'b0}  ;
    assign memory[   77  ] = {16'b0}  ;
    assign memory[   78  ] = {16'b0}  ;
    assign memory[   79  ] = {16'b0}  ;
    assign memory[   80  ] = {16'b0}  ;
    assign memory[   81  ] = {16'b0}  ;
    assign memory[   82  ] = {16'b0}  ;
    assign memory[   83  ] = {16'b0}  ;
    assign memory[   84  ] = {16'b0}  ;
    assign memory[   85  ] = {16'b0}  ;
    assign memory[   86  ] = {16'b0}  ;
    assign memory[   87  ] = {16'b0}  ;
    assign memory[   88  ] = {16'b0}  ;
    assign memory[   89  ] = {16'b0}  ;
    assign memory[   90  ] = {16'b0}  ;
    assign memory[   91  ] = {16'b0}  ;
    assign memory[   92  ] = {16'b0}  ;
    assign memory[   93  ] = {16'b0}  ;
    assign memory[   94  ] = {16'b0}  ;
    assign memory[   95  ] = {16'b0}  ;
    assign memory[   96  ] = {16'b0}  ;
    assign memory[   97  ] = {16'b0}  ;
    assign memory[   98  ] = {16'b0}  ;
    assign memory[   99  ] = {16'b0}  ;
    assign memory[   100  ] = {16'b0}  ;
    assign memory[   101  ] = {16'b0}  ;
    assign memory[   102  ] = {16'b0}  ;
    assign memory[   103  ] = {16'b0}  ;
    assign memory[   104  ] = {16'b0}  ;
    assign memory[   105  ] = {16'b0}  ;
    assign memory[   106  ] = {16'b0}  ;
    assign memory[   107  ] = {16'b0}  ;
    assign memory[   108  ] = {16'b0}  ;
    assign memory[   109  ] = {16'b0}  ;
    assign memory[   110  ] = {16'b0}  ;
    assign memory[   111  ] = {16'b0}  ;
    assign memory[   112  ] = {16'b0}  ;
    assign memory[   113  ] = {16'b0}  ;
    assign memory[   114  ] = {16'b0}  ;
    assign memory[   115  ] = {16'b0}  ;
    assign memory[   116  ] = {16'b0}  ;
    assign memory[   117  ] = {16'b0}  ;
    assign memory[   118  ] = {16'b0}  ;
    assign memory[   119  ] = {16'b0}  ;
    assign memory[   120  ] = {16'b0}  ;
    assign memory[   121  ] = {16'b0}  ;
    assign memory[   122  ] = {16'b0}  ;
    assign memory[   123  ] = {16'b0}  ;
    assign memory[   124  ] = {16'b0}  ;
    assign memory[   125  ] = {16'b0}  ;
    assign memory[   126  ] = {16'b0}  ;
    assign memory[   127  ] = {16'b0}  ;
    assign memory[   128  ] = {16'b0}  ;
    assign memory[   129  ] = {16'b0}  ;
    assign memory[   130  ] = {16'b0}  ;
    assign memory[   131  ] = {16'b0}  ;
    assign memory[   132  ] = {16'b0}  ;
    assign memory[   133  ] = {16'b0}  ;
    assign memory[   134  ] = {16'b0}  ;
    assign memory[   135  ] = {16'b0}  ;
    assign memory[   136  ] = {16'b0}  ;
    assign memory[   137  ] = {16'b0}  ;
    assign memory[   138  ] = {16'b0}  ;
    assign memory[   139  ] = {16'b0}  ;
    assign memory[   140  ] = {16'b0}  ;
    assign memory[   141  ] = {16'b0}  ;
    assign memory[   142  ] = {16'b0}  ;
    assign memory[   143  ] = {16'b0}  ;
    assign memory[   144  ] = {16'b0}  ;
    assign memory[   145  ] = {16'b0}  ;
    assign memory[   146  ] = {16'b0}  ;
    assign memory[   147  ] = {16'b0}  ;
    assign memory[   148  ] = {16'b0}  ;
    assign memory[   149  ] = {16'b0}  ;
    assign memory[   150  ] = {16'b0}  ;
    assign memory[   151  ] = {16'b0}  ;
    assign memory[   152  ] = {16'b0}  ;
    assign memory[   153  ] = {16'b0}  ;
    assign memory[   154  ] = {16'b0}  ;
    assign memory[   155  ] = {16'b0}  ;
    assign memory[   156  ] = {16'b0}  ;
    assign memory[   157  ] = {16'b0}  ;
    assign memory[   158  ] = {16'b0}  ;
    assign memory[   159  ] = {16'b0}  ;
    assign memory[   160  ] = {16'b0}  ;
    assign memory[   161  ] = {16'b0}  ;
    assign memory[   162  ] = {16'b0}  ;
    assign memory[   163  ] = {16'b0}  ;
    assign memory[   164  ] = {16'b0}  ;
    assign memory[   165  ] = {16'b0}  ;
    assign memory[   166  ] = {16'b0}  ;
    assign memory[   167  ] = {16'b0}  ;
    assign memory[   168  ] = {16'b0}  ;
    assign memory[   169  ] = {16'b0}  ;
    assign memory[   170  ] = {16'b0}  ;
    assign memory[   171  ] = {16'b0}  ;
    assign memory[   172  ] = {16'b0}  ;
    assign memory[   173  ] = {16'b0}  ;
    assign memory[   174  ] = {16'b0}  ;
    assign memory[   175  ] = {16'b0}  ;
    assign memory[   176  ] = {16'b0}  ;
    assign memory[   177  ] = {16'b0}  ;
    assign memory[   178  ] = {16'b0}  ;
    assign memory[   179  ] = {16'b0}  ;
    assign memory[   180  ] = {16'b0}  ;
    assign memory[   181  ] = {16'b0}  ;
    assign memory[   182  ] = {16'b0}  ;
    assign memory[   183  ] = {16'b0}  ;
    assign memory[   184  ] = {16'b0}  ;
    assign memory[   185  ] = {16'b0}  ;
    assign memory[   186  ] = {16'b0}  ;
    assign memory[   187  ] = {16'b0}  ;
    assign memory[   188  ] = {16'b0}  ;
    assign memory[   189  ] = {16'b0}  ;
    assign memory[   190  ] = {16'b0}  ;
    assign memory[   191  ] = {16'b0}  ;
    assign memory[   192  ] = {16'b0}  ;
    assign memory[   193  ] = {16'b0}  ;
    assign memory[   194  ] = {16'b0}  ;
    assign memory[   195  ] = {16'b0}  ;
    assign memory[   196  ] = {16'b0}  ;
    assign memory[   197  ] = {16'b0}  ;
    assign memory[   198  ] = {16'b0}  ;
    assign memory[   199  ] = {16'b0}  ;
    assign memory[   200  ] = {16'b0}  ;
    assign memory[   201  ] = {16'b0}  ;
    assign memory[   202  ] = {16'b0}  ;
    assign memory[   203  ] = {16'b0}  ;
    assign memory[   204  ] = {16'b0}  ;
    assign memory[   205  ] = {16'b0}  ;
    assign memory[   206  ] = {16'b0}  ;
    assign memory[   207  ] = {16'b0}  ;
    assign memory[   208  ] = {16'b0}  ;
    assign memory[   209  ] = {16'b0}  ;
    assign memory[   210  ] = {16'b0}  ;
    assign memory[   211  ] = {16'b0}  ;
    assign memory[   212  ] = {16'b0}  ;
    assign memory[   213  ] = {16'b0}  ;
    assign memory[   214  ] = {16'b0}  ;
    assign memory[   215  ] = {16'b0}  ;
    assign memory[   216  ] = {16'b0}  ;
    assign memory[   217  ] = {16'b0}  ;
    assign memory[   218  ] = {16'b0}  ;
    assign memory[   219  ] = {16'b0}  ;
    assign memory[   220  ] = {16'b0}  ;
    assign memory[   221  ] = {16'b0}  ;
    assign memory[   222  ] = {16'b0}  ;
    assign memory[   223  ] = {16'b0}  ;
    assign memory[   224  ] = {16'b0}  ;
    assign memory[   225  ] = {16'b0}  ;
    assign memory[   226  ] = {16'b0}  ;
    assign memory[   227  ] = {16'b0}  ;
    assign memory[   228  ] = {16'b0}  ;
    assign memory[   229  ] = {16'b0}  ;
    assign memory[   230  ] = {16'b0}  ;
    assign memory[   231  ] = {16'b0}  ;
    assign memory[   232  ] = {16'b0}  ;
    assign memory[   233  ] = {16'b0}  ;
    assign memory[   234  ] = {16'b0}  ;
    assign memory[   235  ] = {16'b0}  ;
    assign memory[   236  ] = {16'b0}  ;
    assign memory[   237  ] = {16'b0}  ;
    assign memory[   238  ] = {16'b0}  ;
    assign memory[   239  ] = {16'b0}  ;
    assign memory[   240  ] = {16'b0}  ;
    assign memory[   241  ] = {16'b0}  ;
    assign memory[   242  ] = {16'b0}  ;
    assign memory[   243  ] = {16'b0}  ;
    assign memory[   244  ] = {16'b0}  ;
    assign memory[   245  ] = {16'b0}  ;
    assign memory[   246  ] = {16'b0}  ;
    assign memory[   247  ] = {16'b0}  ;
    assign memory[   248  ] = {16'b0}  ;
    assign memory[   249  ] = {16'b0}  ;
    assign memory[   250  ] = {16'b0}  ;
    assign memory[   251  ] = {16'b0}  ;
    assign memory[   252  ] = {16'b0}  ;
    assign memory[   253  ] = {16'b0}  ;
    assign memory[   254  ] = {16'b0}  ;
    assign memory[   255  ] = {16'b0}  ;
    assign memory[   256  ] = {16'b0}  ;
    assign memory[   257  ] = {16'b0}  ;
    assign memory[   258  ] = {16'b0}  ;
    assign memory[   259  ] = {16'b0}  ;
    assign memory[   260  ] = {16'b0}  ;
    assign memory[   261  ] = {16'b0}  ;
    assign memory[   262  ] = {16'b0}  ;
    assign memory[   263  ] = {16'b0}  ;
    assign memory[   264  ] = {16'b0}  ;
    assign memory[   265  ] = {16'b0}  ;
    assign memory[   266  ] = {16'b0}  ;
    assign memory[   267  ] = {16'b0}  ;
    assign memory[   268  ] = {16'b0}  ;
    assign memory[   269  ] = {16'b0}  ;
    assign memory[   270  ] = {16'b0}  ;
    assign memory[   271  ] = {16'b0}  ;
    assign memory[   272  ] = {16'b0}  ;
    assign memory[   273  ] = {16'b0}  ;
    assign memory[   274  ] = {16'b0}  ;
    assign memory[   275  ] = {16'b0}  ;
    assign memory[   276  ] = {16'b0}  ;
    assign memory[   277  ] = {16'b0}  ;
    assign memory[   278  ] = {16'b0}  ;
    assign memory[   279  ] = {16'b0}  ;
    assign memory[   280  ] = {16'b0}  ;
    assign memory[   281  ] = {16'b0}  ;
    assign memory[   282  ] = {16'b0}  ;
    assign memory[   283  ] = {16'b0}  ;
    assign memory[   284  ] = {16'b0}  ;
    assign memory[   285  ] = {16'b0}  ;
    assign memory[   286  ] = {16'b0}  ;
    assign memory[   287  ] = {16'b0}  ;
    assign memory[   288  ] = {16'b0}  ;
    assign memory[   289  ] = {16'b0}  ;
    assign memory[   290  ] = {16'b0}  ;
    assign memory[   291  ] = {16'b0}  ;
    assign memory[   292  ] = {16'b0}  ;
    assign memory[   293  ] = {16'b0}  ;
    assign memory[   294  ] = {16'b0}  ;
    assign memory[   295  ] = {16'b0}  ;
    assign memory[   296  ] = {16'b0}  ;
    assign memory[   297  ] = {16'b0}  ;
    assign memory[   298  ] = {16'b0}  ;
    assign memory[   299  ] = {16'b0}  ;
    assign memory[   300  ] = {16'b0}  ;
    assign memory[   301  ] = {16'b0}  ;
    assign memory[   302  ] = {16'b0}  ;
    assign memory[   303  ] = {16'b0}  ;
    assign memory[   304  ] = {16'b0}  ;
    assign memory[   305  ] = {16'b0}  ;
    assign memory[   306  ] = {16'b0}  ;
    assign memory[   307  ] = {16'b0}  ;
    assign memory[   308  ] = {16'b0}  ;
    assign memory[   309  ] = {16'b0}  ;
    assign memory[   310  ] = {16'b0}  ;
    assign memory[   311  ] = {16'b0}  ;
    assign memory[   312  ] = {16'b0}  ;
    assign memory[   313  ] = {16'b0}  ;
    assign memory[   314  ] = {16'b0}  ;
    assign memory[   315  ] = {16'b0}  ;
    assign memory[   316  ] = {16'b0}  ;
    assign memory[   317  ] = {16'b0}  ;
    assign memory[   318  ] = {16'b0}  ;
    assign memory[   319  ] = {16'b0}  ;
    assign memory[   320  ] = {16'b0}  ;
    assign memory[   321  ] = {16'b0}  ;
    assign memory[   322  ] = {16'b0}  ;
    assign memory[   323  ] = {16'b0}  ;
    assign memory[   324  ] = {16'b0}  ;
    assign memory[   325  ] = {16'b0}  ;
    assign memory[   326  ] = {16'b0}  ;
    assign memory[   327  ] = {16'b0}  ;
    assign memory[   328  ] = {16'b0}  ;
    assign memory[   329  ] = {16'b0}  ;
    assign memory[   330  ] = {16'b0}  ;
    assign memory[   331  ] = {16'b0}  ;
    assign memory[   332  ] = {16'b0}  ;
    assign memory[   333  ] = {16'b0}  ;
    assign memory[   334  ] = {16'b0}  ;
    assign memory[   335  ] = {16'b0}  ;
    assign memory[   336  ] = {16'b0}  ;
    assign memory[   337  ] = {16'b0}  ;
    assign memory[   338  ] = {16'b0}  ;
    assign memory[   339  ] = {16'b0}  ;
    assign memory[   340  ] = {16'b0}  ;
    assign memory[   341  ] = {16'b0}  ;
    assign memory[   342  ] = {16'b0}  ;
    assign memory[   343  ] = {16'b0}  ;
    assign memory[   344  ] = {16'b0}  ;
    assign memory[   345  ] = {16'b0}  ;
    assign memory[   346  ] = {16'b0}  ;
    assign memory[   347  ] = {16'b0}  ;
    assign memory[   348  ] = {16'b0}  ;
    assign memory[   349  ] = {16'b0}  ;
    assign memory[   350  ] = {16'b0}  ;
    assign memory[   351  ] = {16'b0}  ;
    assign memory[   352  ] = {16'b0}  ;
    assign memory[   353  ] = {16'b0}  ;
    assign memory[   354  ] = {16'b0}  ;
    assign memory[   355  ] = {16'b0}  ;
    assign memory[   356  ] = {16'b0}  ;
    assign memory[   357  ] = {16'b0}  ;
    assign memory[   358  ] = {16'b0}  ;
    assign memory[   359  ] = {16'b0}  ;
    assign memory[   360  ] = {16'b0}  ;
    assign memory[   361  ] = {16'b0}  ;
    assign memory[   362  ] = {16'b0}  ;
    assign memory[   363  ] = {16'b0}  ;
    assign memory[   364  ] = {16'b0}  ;
    assign memory[   365  ] = {16'b0}  ;
    assign memory[   366  ] = {16'b0}  ;
    assign memory[   367  ] = {16'b0}  ;
    assign memory[   368  ] = {16'b0}  ;
    assign memory[   369  ] = {16'b0}  ;
    assign memory[   370  ] = {16'b0}  ;
    assign memory[   371  ] = {16'b0}  ;
    assign memory[   372  ] = {16'b0}  ;
    assign memory[   373  ] = {16'b0}  ;
    assign memory[   374  ] = {16'b0}  ;
    assign memory[   375  ] = {16'b0}  ;
    assign memory[   376  ] = {16'b0}  ;
    assign memory[   377  ] = {16'b0}  ;
    assign memory[   378  ] = {16'b0}  ;
    assign memory[   379  ] = {16'b0}  ;
    assign memory[   380  ] = {16'b0}  ;
    assign memory[   381  ] = {16'b0}  ;
    assign memory[   382  ] = {16'b0}  ;
    assign memory[   383  ] = {16'b0}  ;
    assign memory[   384  ] = {16'b0}  ;
    assign memory[   385  ] = {16'b0}  ;
    assign memory[   386  ] = {16'b0}  ;
    assign memory[   387  ] = {16'b0}  ;
    assign memory[   388  ] = {16'b0}  ;
    assign memory[   389  ] = {16'b0}  ;
    assign memory[   390  ] = {16'b0}  ;
    assign memory[   391  ] = {16'b0}  ;
    assign memory[   392  ] = {16'b0}  ;
    assign memory[   393  ] = {16'b0}  ;
    assign memory[   394  ] = {16'b0}  ;
    assign memory[   395  ] = {16'b0}  ;
    assign memory[   396  ] = {16'b0}  ;
    assign memory[   397  ] = {16'b0}  ;
    assign memory[   398  ] = {16'b0}  ;
    assign memory[   399  ] = {16'b0}  ;
    assign memory[   400  ] = {16'b0}  ;
    assign memory[   401  ] = {16'b0}  ;
    assign memory[   402  ] = {16'b0}  ;
    assign memory[   403  ] = {16'b0}  ;
    assign memory[   404  ] = {16'b0}  ;
    assign memory[   405  ] = {16'b0}  ;
    assign memory[   406  ] = {16'b0}  ;
    assign memory[   407  ] = {16'b0}  ;
    assign memory[   408  ] = {16'b0}  ;
    assign memory[   409  ] = {16'b0}  ;
    assign memory[   410  ] = {16'b0}  ;
    assign memory[   411  ] = {16'b0}  ;
    assign memory[   412  ] = {16'b0}  ;
    assign memory[   413  ] = {16'b0}  ;
    assign memory[   414  ] = {16'b0}  ;
    assign memory[   415  ] = {16'b0}  ;
    assign memory[   416  ] = {16'b0}  ;
    assign memory[   417  ] = {16'b0}  ;
    assign memory[   418  ] = {16'b0}  ;
    assign memory[   419  ] = {16'b0}  ;
    assign memory[   420  ] = {16'b0}  ;
    assign memory[   421  ] = {16'b0}  ;
    assign memory[   422  ] = {16'b0}  ;
    assign memory[   423  ] = {16'b0}  ;
    assign memory[   424  ] = {16'b0}  ;
    assign memory[   425  ] = {16'b0}  ;
    assign memory[   426  ] = {16'b0}  ;
    assign memory[   427  ] = {16'b0}  ;
    assign memory[   428  ] = {16'b0}  ;
    assign memory[   429  ] = {16'b0}  ;
    assign memory[   430  ] = {16'b0}  ;
    assign memory[   431  ] = {16'b0}  ;
    assign memory[   432  ] = {16'b0}  ;
    assign memory[   433  ] = {16'b0}  ;
    assign memory[   434  ] = {16'b0}  ;
    assign memory[   435  ] = {16'b0}  ;
    assign memory[   436  ] = {16'b0}  ;
    assign memory[   437  ] = {16'b0}  ;
    assign memory[   438  ] = {16'b0}  ;
    assign memory[   439  ] = {16'b0}  ;
    assign memory[   440  ] = {16'b0}  ;
    assign memory[   441  ] = {16'b0}  ;
    assign memory[   442  ] = {16'b0}  ;
    assign memory[   443  ] = {16'b0}  ;
    assign memory[   444  ] = {16'b0}  ;
    assign memory[   445  ] = {16'b0}  ;
    assign memory[   446  ] = {16'b0}  ;
    assign memory[   447  ] = {16'b0}  ;
    assign memory[   448  ] = {16'b0}  ;
    assign memory[   449  ] = {16'b0}  ;
    assign memory[   450  ] = {16'b0}  ;
    assign memory[   451  ] = {16'b0}  ;
    assign memory[   452  ] = {16'b0}  ;
    assign memory[   453  ] = {16'b0}  ;
    assign memory[   454  ] = {16'b0}  ;
    assign memory[   455  ] = {16'b0}  ;
    assign memory[   456  ] = {16'b0}  ;
    assign memory[   457  ] = {16'b0}  ;
    assign memory[   458  ] = {16'b0}  ;
    assign memory[   459  ] = {16'b0}  ;
    assign memory[   460  ] = {16'b0}  ;
    assign memory[   461  ] = {16'b0}  ;
    assign memory[   462  ] = {16'b0}  ;
    assign memory[   463  ] = {16'b0}  ;
    assign memory[   464  ] = {16'b0}  ;
    assign memory[   465  ] = {16'b0}  ;
    assign memory[   466  ] = {16'b0}  ;
    assign memory[   467  ] = {16'b0}  ;
    assign memory[   468  ] = {16'b0}  ;
    assign memory[   469  ] = {16'b0}  ;
    assign memory[   470  ] = {16'b0}  ;
    assign memory[   471  ] = {16'b0}  ;
    assign memory[   472  ] = {16'b0}  ;
    assign memory[   473  ] = {16'b0}  ;
    assign memory[   474  ] = {16'b0}  ;
    assign memory[   475  ] = {16'b0}  ;
    assign memory[   476  ] = {16'b0}  ;
    assign memory[   477  ] = {16'b0}  ;
    assign memory[   478  ] = {16'b0}  ;
    assign memory[   479  ] = {16'b0}  ;
    assign memory[   480  ] = {16'b0}  ;
    assign memory[   481  ] = {16'b0}  ;
    assign memory[   482  ] = {16'b0}  ;
    assign memory[   483  ] = {16'b0}  ;
    assign memory[   484  ] = {16'b0}  ;
    assign memory[   485  ] = {16'b0}  ;
    assign memory[   486  ] = {16'b0}  ;
    assign memory[   487  ] = {16'b0}  ;
    assign memory[   488  ] = {16'b0}  ;
    assign memory[   489  ] = {16'b0}  ;
    assign memory[   490  ] = {16'b0}  ;
    assign memory[   491  ] = {16'b0}  ;
    assign memory[   492  ] = {16'b0}  ;
    assign memory[   493  ] = {16'b0}  ;
    assign memory[   494  ] = {16'b0}  ;
    assign memory[   495  ] = {16'b0}  ;
    assign memory[   496  ] = {16'b0}  ;
    assign memory[   497  ] = {16'b0}  ;
    assign memory[   498  ] = {16'b0}  ;
    assign memory[   499  ] = {16'b0}  ;
    assign memory[   500  ] = {16'b0}  ;
    assign memory[   501  ] = {16'b0}  ;
    assign memory[   502  ] = {16'b0}  ;
    assign memory[   503  ] = {16'b0}  ;
    assign memory[   504  ] = {16'b0}  ;
    assign memory[   505  ] = {16'b0}  ;
    assign memory[   506  ] = {16'b0}  ;
    assign memory[   507  ] = {16'b0}  ;
    assign memory[   508  ] = {16'b0}  ;
    assign memory[   509  ] = {16'b0}  ;
    assign memory[   510  ] = {16'b0}  ;
    assign memory[   511  ] = {16'b0}  ;

endmodule       
